library verilog;
use verilog.vl_types.all;
entity project_tb is
end project_tb;
