library verilog;
use verilog.vl_types.all;
entity tap_tb is
end tap_tb;
